//define key codes
`define KEY_1 4'd1
`define KEY_2 4'd2
`define KEY_3 4'd3
`define KEY_4 4'd4
`define KEY_5 4'd5
`define KEY_6 4'd6
`define KEY_7 4'd7
`define KEY_8 4'd8
`define KEY_9 4'd9
`define KEY_0 4'd0
`define KEY_ADD 4'd11
`define KEY_SUBTRACT 4'd12
`define KEY_MULTIPLY 4'd13
`define KEY_ENTER 4'd14
`define KEY_CLEAR 4'd15

//define state code
`define STAT_DIGIT3 3'd0
`define STAT_DIGIT2 3'd1
`define STAT_OPERATOR 3'd2
`define STAT_DIGIT1 3'd3
`define STAT_DIGIT0 3'd4
`define STAT_DISPLAY 3'd5


